module mult256(in,out);
	input [31:0] in;
	output [31:0] out;
	assign out = in * 32'd256;
endmodule