// Copyright (C) 1991-2009 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 9.0 Build 132 02/25/2009 SJ Full Version
// Created on Sat Dec 29 12:57:10 2012

// synthesis message_off 10175

`timescale 1ns/1ns

module SM1 (
    reset,clock,start,usedw1a32,empty1a,nioswrite,empty3Re,empty2Re,empty5,empty4a,full4a,full4b,full5,usedw1b64,f642Re,usedw1a64,usedw2Re64,usedw3Re64,
    wrreq1a,wrreq1b,rdreq1a,rdreq1b,wrreq2,niosread2,rdreq3,wrreq4a,wrreq4b,rdreq4,wrreq5,niosread5,fft_enable,selmuxFIFO,selmuxFFT);

    input reset;
    input clock;
    input start;
    input usedw1a32;
    input empty1a;
    input nioswrite;
    input empty3Re;
    input empty2Re;
    input empty5;
    input empty4a;
    input full4a;
    input full4b;
    input full5;
    input usedw1b64;
    input f642Re;
    input usedw1a64;
    input usedw2Re64;
    input usedw3Re64;
    tri0 reset;
    tri0 start;
    tri0 usedw1a32;
    tri0 empty1a;
    tri0 nioswrite;
    tri0 empty3Re;
    tri0 empty2Re;
    tri0 empty5;
    tri0 empty4a;
    tri0 full4a;
    tri0 full4b;
    tri0 full5;
    tri0 usedw1b64;
    tri0 f642Re;
    tri0 usedw1a64;
    tri0 usedw2Re64;
    tri0 usedw3Re64;
    output wrreq1a;
    output wrreq1b;
    output rdreq1a;
    output rdreq1b;
    output wrreq2;
    output niosread2;
    output rdreq3;
    output wrreq4a;
    output wrreq4b;
    output rdreq4;
    output wrreq5;
    output niosread5;
    output fft_enable;
    output selmuxFIFO;
    output selmuxFFT;
    reg wrreq1a;
    reg wrreq1b;
    reg rdreq1a;
    reg reg_rdreq1a;
    reg rdreq1b;
    reg reg_rdreq1b;
    reg wrreq2;
    reg reg_wrreq2;
    reg niosread2;
    reg reg_niosread2;
    reg rdreq3;
    reg reg_rdreq3;
    reg wrreq4a;
    reg reg_wrreq4a;
    reg wrreq4b;
    reg reg_wrreq4b;
    reg rdreq4;
    reg reg_rdreq4;
    reg wrreq5;
    reg reg_wrreq5;
    reg niosread5;
    reg reg_niosread5;
    reg fft_enable;
    reg reg_fft_enable;
    reg selmuxFIFO;
    reg reg_selmuxFIFO;
    reg selmuxFFT;
    reg reg_selmuxFFT;
    reg [15:0] fstate;
    reg [15:0] reg_fstate;
    parameter idle=0,S1=1,S2=2,S3=3,S4=4,S5=5,S6=6,S7=7,S8=8,S9=9,S10=10,S11=11,S12=12,S13=13,S14=14,S1_1=15;

    initial
    begin
        reg_rdreq1a <= 1'b0;
        reg_rdreq1b <= 1'b0;
        reg_wrreq2 <= 1'b0;
        reg_niosread2 <= 1'b0;
        reg_rdreq3 <= 1'b0;
        reg_wrreq4a <= 1'b0;
        reg_wrreq4b <= 1'b0;
        reg_rdreq4 <= 1'b0;
        reg_wrreq5 <= 1'b0;
        reg_niosread5 <= 1'b0;
        reg_fft_enable <= 1'b0;
        reg_selmuxFIFO <= 1'b0;
        reg_selmuxFFT <= 1'b0;
    end

    always @(posedge clock or negedge reset)
    begin
        if (~reset) begin
            fstate <= idle;
        end
        else begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or start or usedw1a32 or empty1a or nioswrite or empty3Re or empty2Re or empty5 or empty4a or full4a or full4b or full5 or usedw1b64 or f642Re or usedw1a64 or usedw2Re64 or usedw3Re64 or reg_rdreq1a or reg_rdreq1b or reg_wrreq2 or reg_niosread2 or reg_rdreq3 or reg_wrreq4a or reg_wrreq4b or reg_rdreq4 or reg_wrreq5 or reg_niosread5 or reg_fft_enable or reg_selmuxFIFO or reg_selmuxFFT)
    begin
        wrreq1a <= 1'b0;
        wrreq1b <= 1'b0;
        reg_rdreq1a <= 1'b0;
        reg_rdreq1b <= 1'b0;
        reg_wrreq2 <= 1'b0;
        reg_niosread2 <= 1'b0;
        reg_rdreq3 <= 1'b0;
        reg_wrreq4a <= 1'b0;
        reg_wrreq4b <= 1'b0;
        reg_rdreq4 <= 1'b0;
        reg_wrreq5 <= 1'b0;
        reg_niosread5 <= 1'b0;
        reg_fft_enable <= 1'b0;
        reg_selmuxFIFO <= 1'b0;
        reg_selmuxFFT <= 1'b0;
        rdreq1a <= 1'b0;
        rdreq1b <= 1'b0;
        wrreq2 <= 1'b0;
        niosread2 <= 1'b0;
        rdreq3 <= 1'b0;
        wrreq4a <= 1'b0;
        wrreq4b <= 1'b0;
        rdreq4 <= 1'b0;
        wrreq5 <= 1'b0;
        niosread5 <= 1'b0;
        fft_enable <= 1'b0;
        selmuxFIFO <= 1'b0;
        selmuxFFT <= 1'b0;
        case (fstate)
            idle: begin
                if ((start == 1'b1))
                    reg_fstate <= S1;
                else if ((start == 1'b0))
                    reg_fstate <= idle;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= idle;

                wrreq1a <= 1'b0;

                wrreq1b <= 1'b0;

                reg_rdreq1a <= 1'b0;

                reg_rdreq1b <= 1'b0;

                reg_wrreq2 <= 1'b0;

                reg_niosread2 <= 1'b0;

                reg_rdreq3 <= 1'b0;

                reg_wrreq4a <= 1'b0;

                reg_wrreq4b <= 1'b0;

                reg_rdreq4 <= 1'b0;

                reg_wrreq5 <= 1'b0;

                reg_niosread5 <= 1'b0;

                reg_fft_enable <= 1'b0;

                reg_selmuxFIFO <= 1'b0;

                reg_selmuxFFT <= 1'b0;
            end
            S1: begin
                if ((usedw1a32 == 1'b0))
                    reg_fstate <= S1;
                else if ((usedw1a32 == 1'b1))
                    reg_fstate <= S1_1;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= S1;

                wrreq1a <= 1'b1;

                if ((usedw1a32 == 1'b1))
                    wrreq1b <= 1'b1;
                // Inserting 'else' block to prevent latch inference
                else
                    wrreq1b <= 1'b0;
            end
            S2: begin
                if ((empty1a == 1'b1))
                    reg_fstate <= S3;
                else if ((empty1a == 1'b0))
                    reg_fstate <= S2;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= S2;

                if ((usedw1b64 == 1'b0))
                    wrreq1b <= 1'b1;
                // Inserting 'else' block to prevent latch inference
                else
                    wrreq1b <= 1'b0;

                reg_rdreq1a <= 1'b1;

                reg_fft_enable <= 1'b1;
            end
            S3: begin
                if ((usedw2Re64 == 1'b1))
                    reg_fstate <= S4;
                else if ((usedw2Re64 == 1'b0))
                    reg_fstate <= S3;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= S3;

                if ((usedw1b64 == 1'b1))
                    wrreq1b <= 1'b0;
                // Inserting 'else' block to prevent latch inference
                else
                    wrreq1b <= 1'b0;

                reg_rdreq1a <= 1'b0;

                reg_rdreq1b <= 1'b1;

                reg_wrreq2 <= 1'b1;

                reg_fft_enable <= 1'b1;

                reg_selmuxFIFO <= 1'b1;
            end
            S4: begin
                if ((f642Re == 1'b1))
                    reg_fstate <= S5;
                else if ((f642Re == 1'b0))
                    reg_fstate <= S4;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= S4;

                reg_rdreq1b <= 1'b0;

                reg_wrreq2 <= 1'b1;

                reg_niosread2 <= 1'b1;

                reg_fft_enable <= 1'b0;
            end
            S5: begin
                if ((empty2Re == 1'b1))
                    reg_fstate <= S6;
                else if ((empty2Re == 1'b0))
                    reg_fstate <= S5;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= S5;

                reg_wrreq2 <= 1'b0;

                reg_niosread2 <= 1'b1;
            end
            S6: begin
                if ((nioswrite == 1'b0))
                    reg_fstate <= S6;
                else if ((nioswrite == 1'b1))
                    reg_fstate <= S7;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= S6;

                reg_niosread2 <= 1'b0;

                reg_selmuxFIFO <= 1'b0;
            end
            S7: begin
                if ((usedw3Re64 == 1'b0))
                    reg_fstate <= S7;
                else if ((usedw3Re64 == 1'b1))
                    reg_fstate <= S8;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= S7;

                reg_selmuxFFT <= 1'b1;
            end
            S8: begin
                if ((empty3Re == 1'b0))
                    reg_fstate <= S8;
                else if ((empty3Re == 1'b1))
                    reg_fstate <= S9;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= S8;

                reg_rdreq3 <= 1'b1;

                reg_fft_enable <= 1'b1;

                reg_selmuxFFT <= 1'b1;
            end
            S9: begin
                if ((full4a == 1'b0))
                    reg_fstate <= S9;
                else if ((full4a == 1'b1))
                    reg_fstate <= S10;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= S9;

                reg_wrreq4a <= 1'b1;

                reg_selmuxFFT <= 1'b1;
            end
            S10: begin
                if ((full4b == 1'b0))
                    reg_fstate <= S10;
                else if ((full4b == 1'b1))
                    reg_fstate <= S11;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= S10;

                reg_wrreq4a <= 1'b0;

                reg_wrreq4b <= 1'b1;

                reg_selmuxFIFO <= 1'b1;

                reg_selmuxFFT <= 1'b1;
            end
            S11: begin
                if ((empty4a == 1'b0))
                    reg_fstate <= S11;
                else if ((empty4a == 1'b1))
                    reg_fstate <= S12;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= S11;

                reg_rdreq4 <= 1'b1;

                reg_selmuxFIFO <= 1'b0;

                reg_selmuxFFT <= 1'b1;
            end
            S12: begin
                if ((full5 == 1'b1))
                    reg_fstate <= S13;
                else if ((full5 == 1'b0))
                    reg_fstate <= S12;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= S12;

                reg_rdreq4 <= 1'b0;

                reg_wrreq5 <= 1'b1;
            end
            S13: begin
                if ((empty5 == 1'b1))
                    reg_fstate <= S14;
                else if ((empty5 == 1'b0))
                    reg_fstate <= S13;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= S13;

                reg_wrreq5 <= 1'b0;

                reg_niosread5 <= 1'b1;
            end
            S14: begin
                if ((start == 1'b1))
                    reg_fstate <= S1;
                else if ((start == 1'b0))
                    reg_fstate <= S14;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= S14;

                reg_niosread5 <= 1'b0;

                reg_fft_enable <= 1'b0;

                reg_selmuxFFT <= 1'b0;
            end
            S1_1: begin
                if ((usedw1a64 == 1'b1))
                    reg_fstate <= S2;
                else if ((usedw1a64 == 1'b0))
                    reg_fstate <= S1_1;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= S1_1;

                wrreq1a <= 1'b1;

                wrreq1b <= 1'b1;
            end
            default: begin
                wrreq1a <= 1'bx;
                wrreq1b <= 1'bx;
                reg_rdreq1a <= 1'bx;
                reg_rdreq1b <= 1'bx;
                reg_wrreq2 <= 1'bx;
                reg_niosread2 <= 1'bx;
                reg_rdreq3 <= 1'bx;
                reg_wrreq4a <= 1'bx;
                reg_wrreq4b <= 1'bx;
                reg_rdreq4 <= 1'bx;
                reg_wrreq5 <= 1'bx;
                reg_niosread5 <= 1'bx;
                reg_fft_enable <= 1'bx;
                reg_selmuxFIFO <= 1'bx;
                reg_selmuxFFT <= 1'bx;
                $display ("Reach undefined state");
            end
        endcase
        rdreq1a <= reg_rdreq1a;
        rdreq1b <= reg_rdreq1b;
        wrreq2 <= reg_wrreq2;
        niosread2 <= reg_niosread2;
        rdreq3 <= reg_rdreq3;
        wrreq4a <= reg_wrreq4a;
        wrreq4b <= reg_wrreq4b;
        rdreq4 <= reg_rdreq4;
        wrreq5 <= reg_wrreq5;
        niosread5 <= reg_niosread5;
        fft_enable <= reg_fft_enable;
        selmuxFIFO <= reg_selmuxFIFO;
        selmuxFFT <= reg_selmuxFFT;
    end
endmodule // SM1
